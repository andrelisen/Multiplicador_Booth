library verilog;
use verilog.vl_types.all;
entity Mult_Booth_PC_vlg_vec_tst is
end Mult_Booth_PC_vlg_vec_tst;
