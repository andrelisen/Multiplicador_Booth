library verilog;
use verilog.vl_types.all;
entity Mult_Booth_PO_vlg_vec_tst is
end Mult_Booth_PO_vlg_vec_tst;
